`timescale 1ns/1ps

// =============================================================================
// Module: TimeSurfaceBinning
// =============================================================================
// Spatio-Temporal Pooling for DVS Gesture Classification
//
// Description:
//   Accumulates DVS events into a ring buffer of 2D histograms (bins) over time.
//   Periodically rotates bins based on timestamps.
//   Flattens the most recent N bins into a vector for classification.
//
// Parameters:
//   CLK_FREQ_HZ     - System clock frequency
//   WINDOW_MS       - Total duration of the observation window (e.g., 400ms)
//   NUM_BINS        - Number of bins in the ring buffer (e.g., 8)
//   READOUT_BINS    - Number of bins to read out for classification (e.g., 5)
//                     Must be <= NUM_BINS.
//   GRID_SIZE       - Spatial grid dimension (e.g., 16x16)
//   COUNTER_BITS    - Bit width for event counters in each bin cell
//
// =============================================================================

module TimeSurfaceBinning #(
    parameter CLK_FREQ_HZ     = 12_000_000,
    parameter WINDOW_MS       = 400,
    parameter NUM_BINS        = 8,
    parameter READOUT_BINS    = 5,
    parameter GRID_SIZE       = 16,
    parameter COUNTER_BITS    = 8
)(
    input  logic        clk,
    input  logic        rst,

    // Input DVS Events (from SpatialCompressor)
    input  logic        event_valid,
    input  logic signed [4:0] event_x,   // [-8 to +7] relative to center
    input  logic signed [4:0] event_y,   // [-8 to +7] relative to center
    input  logic        event_polarity,

    // Timing Logic (using internal cycle counter for simplicity, approximating timestamps)
    // In a real system, we might use the event timestamp, but here we count cycles
    // to determine bin boundaries as per the param description "window W is split into identical, sequential bins".
    
    // Output to Systolic Array
    // Interface matches the 'feature_in' stream expectation of the systolic array
    output logic        readout_start,              // Pulse to start systolic array
    output logic [COUNTER_BITS-1:0] readout_data,   // Streamed feature data
    output logic        readout_valid               // Data valid qualifier
);

    // =========================================================================
    // Parameters & Derived Constants
    // =========================================================================
    localparam integer BIN_DURATION_MS = WINDOW_MS / NUM_BINS;
    localparam integer CYCLES_PER_BIN  = (CLK_FREQ_HZ / 1000) * BIN_DURATION_MS;
    localparam integer TIMER_BITS      = $clog2(CYCLES_PER_BIN + 1);
    
    localparam integer CELLS_PER_BIN   = GRID_SIZE * GRID_SIZE;
    localparam integer TOTAL_CELLS     = NUM_BINS * CELLS_PER_BIN;
    localparam integer CELL_ADDR_BITS  = $clog2(TOTAL_CELLS);
    localparam integer BIN_IDX_BITS    = $clog2(NUM_BINS);
    localparam integer GRID_ADDR_BITS  = $clog2(CELLS_PER_BIN);

    // =========================================================================
    // Bin Timing & Management
    // =========================================================================
    logic [TIMER_BITS-1:0]   bin_timer;
    logic [BIN_IDX_BITS-1:0] current_bin_idx;  // The bin currently being filled (head)
    
    // Ring Buffer RAM
    // We need to read/modify/write for event accumulation
    // We need to read for readout (potentially concurrent, but we can serialize)
    // Structure: Simple Dual Port RAM (Read and write ports) or just register array if small enough?
    // Total bits = 8 bins * 256 cells * 8 bits = 16Kb. Fits in BRAM.
    // However, simultaneous access might be tricky if an event comes during readout.
    // Priority: Event accumulation has priority to avoid dropping events? 
    // Or Readout has priority?
    // Let's use a standard construct.
    
    logic [COUNTER_BITS-1:0] mem [0:TOTAL_CELLS-1]; // Inferred RAM
    
    // Event Processing Signals
    logic [BIN_IDX_BITS-1:0] event_bin_idx;
    logic [3:0]              mapped_x, mapped_y; // Unsigned [0-15]
    logic [GRID_ADDR_BITS-1:0] event_cell_addr;
    logic [CELL_ADDR_BITS-1:0] event_full_addr;
    
    // Coordinate mapping: input is [-8, +7], center at 0.
    // Map to [0, 15] for indexing.
    // -8 -> 0, +7 -> 15. Add 8.
    assign mapped_x = event_x + 5'd8;
    assign mapped_y = event_y + 5'd8;
    assign event_cell_addr = {mapped_y[3:0], mapped_x[3:0]}; // y*16 + x
    
    // Readout State Machine Signals
    typedef enum logic [1:0] {
        S_IDLE,
        S_READOUT,
        S_CLEAR // We need to clear old bins?
                // Actually, the prompt says "When a bin is filled... clear appropriate memory"
                // Efficient way: clear the *next* bin in the ring before we start filling it?
                // Or clear it as we step into it.
                // Let's implement a clear state that runs when we switch bins.
    } state_t;
    
    state_t state;
    
    // Readout Counters
    logic [BIN_IDX_BITS-1:0] readout_bin_ptr; // Logical bin index (0 to READOUT_BINS-1)
    logic [GRID_ADDR_BITS-1:0] readout_cell_ctr;
    
    // Clear Counters
    logic [GRID_ADDR_BITS-1:0] clear_cell_ctr;
    
    // Flag to trigger readout
    logic trigger_readout;
    
    // =========================================================================
    // Bin Rotation Timer
    // =========================================================================
    always_ff @(posedge clk) begin
        if (rst) begin
            bin_timer <= '0;
            current_bin_idx <= '0;
            trigger_readout <= 1'b0;
            state <= S_CLEAR; // Start by clearing the first bin (or all)
            clear_cell_ctr <= '0;
        end else begin
            trigger_readout <= 1'b0; // Default
            
            // State Machine for Timer / Bin Management
            if (state == S_IDLE || state == S_READOUT) begin
                if (bin_timer >= CYCLES_PER_BIN - 1) begin
                    bin_timer <= '0;
                    
                    // Move to next bin
                    if (current_bin_idx == NUM_BINS - 1)
                        current_bin_idx <= '0;
                    else
                        current_bin_idx <= current_bin_idx + 1'b1;
                        
                    // Check if we have enough history to readout
                    // Prompt says: "When a bin is filled... window W will be matrix covering last B bins"
                    // "If there are not 5 bins in memory yet, skip producing"
                    // For simplicity, we assume valid after initial fill or just always output (zeros effectively).
                    // We trigger readout on every bin switch.
                    trigger_readout <= 1'b1;
                    
                    // We need to clear the NEW bin we just entered to ensure it's fresh for new events
                    // So we transition to a CLEAR state or handle it.
                    // To avoid blocking events for too long, we could clear it "lazy" or use a VALID bit?
                    // RAM method requires write cycles.
                    // Let's use a state to clear it fast. 256 cycles. 
                    // 256 cycles at 12Mhz is ~21us. Bin is ~50ms. Negligible dead time?
                    // Maybe. Let's do it.
                    state <= S_CLEAR;
                    clear_cell_ctr <= '0;
                end else begin
                    bin_timer <= bin_timer + 1'b1;
                end
            end else if (state == S_CLEAR) begin
                // In clear state, we hold the timer? Or keep counting?
                // Probably keep counting to keep real-time accuracy, but if clear phase is short it's fine.
                // Let's pause timer to avoid complexity, error is small.
                if (clear_cell_ctr == CELLS_PER_BIN - 1) begin
                    state <= S_IDLE; // Done clearing
                    // Note: If readout was triggered, we might want to go to READOUT?
                    // But Readout and Clear can happen somewhat in parallel or sequence.
                    // Let's assume Readout is handled by a separate process or interleaved.
                    // To simplify: Main FSM handles Clearing (blocking writes).
                    // Readout FSM handles Reading (reads).
                    // Single port RAM -> Contention.
                    // We really need dual port here if we want to read while writing.
                    // For this exercise, let's assume we can share or block.
                    // "Event comes in... timestamp checked"
                end
                clear_cell_ctr <= clear_cell_ctr + 1'b1;
            end
        end
    end

    // =========================================================================
    // Memory & R/W Logic
    // =========================================================================
    
    // We need to handle:
    // 1. Event Write (Read-Modify-Write increment)
    // 2. Clear Write (Write 0)
    // 3. Readout Read (Read)
    
    // Prioritize: Clear > Event > Readout?
    // Actually, Clear is critical when switching bins.
    
    logic ram_wen;
    logic [CELL_ADDR_BITS-1:0] ram_addr;
    logic [COUNTER_BITS-1:0] ram_wdata;
    logic [COUNTER_BITS-1:0] ram_rdata;
    
    // Logic for pointers
    // Readout of "Last 5 bins".
    // If current_bin_idx is 3. We want bins [3, 2, 1, 0, 7] (most recent first? or chronological?)
    // "flattened... covering the last B bins"
    // Usually chronological: [Oldest ... Newest].
    // Newest is the one just finished? Or the one being filled?
    // "When a bin is filled... last B bins" -> Includes the one just filled.
    // So if we just finished bin 3.
    // Sequence: Bin 7 (Old), Bin 0, Bin 1, Bin 2, Bin 3 (New).
    
    // Readout State Machine
    logic readout_busy;
    logic [BIN_IDX_BITS-1:0] rd_bin_offset; // 0 to READOUT_BINS-1
    logic [GRID_ADDR_BITS-1:0] rd_cell_ctr;
    
    always_ff @(posedge clk) begin
        if (rst) begin
            readout_busy <= 1'b0;
            readout_start <= 1'b0;
            rd_bin_offset <= '0;
            rd_cell_ctr <= '0;
        end else begin
            readout_start <= 1'b0;

            if (trigger_readout) begin
                readout_busy <= 1'b1;
                readout_start <= 1'b1; // Signal start of stream
                rd_bin_offset <= '0;
                rd_cell_ctr <= '0;
            end else if (readout_busy) begin
                // Advance counters (readout_valid driven by assign from readout_valid_d)
                if (rd_cell_ctr == CELLS_PER_BIN - 1) begin
                    rd_cell_ctr <= '0;
                    if (rd_bin_offset == READOUT_BINS - 1) begin
                        readout_busy <= 1'b0;
                    end else begin
                        rd_bin_offset <= rd_bin_offset + 1'b1;
                    end
                end else begin
                    rd_cell_ctr <= rd_cell_ctr + 1'b1;
                end
            end
        end
    end
    
    // Readout Address Calculation
    // We want the OLDEST bin first? Or NEWEST?
    // Matrix usually [Time, Space].
    // Let's assume chronological order [T-4, T-3, T-2, T-1, T-0]
    // T-0 is the bin just completed.
    // current_bin_idx is the *new* empty bin we just switched to.
    // So T-0 is (current_bin_idx - 1).
    // Start bin = (current_bin_idx - 1) - (READOUT_BINS - 1) = current - READOUT_BINS.
    
    // To handle wrap around logic properly:
    // virtual_idx = current_bin_idx + NUM_BINS - READOUT_BINS + rd_bin_offset;
    // actual_idx = virtual_idx % NUM_BINS;
    
    logic [BIN_IDX_BITS:0] calc_bin_idx; // Extra bit for overflow
    logic [BIN_IDX_BITS-1:0] actual_rd_bin_idx;
    
    always_comb begin
        // The bin we just finished filling is (current_bin_idx - 1) modulo NUM_BINS.
        // We want to start reading from (current_bin_idx - READOUT_BINS).
        // Example: N=8, R=5. Cur=2 (just started). Finished=1.
        // We want bins: 5, 6, 7, 0, 1.
        // 2 + 8 - 5 = 5. Offset 0 -> 5. Offset 4 -> 9%8=1. Correct.
        calc_bin_idx = current_bin_idx + NUM_BINS - READOUT_BINS + rd_bin_offset;
        if (calc_bin_idx >= NUM_BINS) 
            actual_rd_bin_idx = calc_bin_idx - NUM_BINS;
        else 
            actual_rd_bin_idx = calc_bin_idx[BIN_IDX_BITS-1:0];
    end

    // RAM Access Arbitration & Address Muxing
    // RAM latency is 1 cycle for read.
    // We need `readout_data` assigned from `mem[addr]`.
    
    // Event Access Logic
    // We need to Read-Modify-Write. This takes 2 cycles for single port RAM.
    // Or we rely on the fact that events are sparse?
    // If we use dual port RAM:
    // Port A: Read/Write for Events/Clearing.
    // Port B: Read for Readout.
    // This allows Readout to happen in parallel with Event integration.
    // However, Clearing (State S_CLEAR) needs to write.
    
    // Let's infer a simple memory block and handle assignments explicitly
    logic [CELL_ADDR_BITS-1:0] clear_addr;
    logic [CELL_ADDR_BITS-1:0] evt_addr; 
    logic [CELL_ADDR_BITS-1:0] rd_addr;
    
    assign clear_addr = {current_bin_idx, clear_cell_ctr};
    assign evt_addr   = {current_bin_idx, event_cell_addr};
    assign rd_addr    = {actual_rd_bin_idx, rd_cell_ctr};

    // Output assignments
    assign readout_data = ram_rdata; // Latched from RAM
    
    // =========================================================================
    // Dual-Port BRAM Implementation
    // Port A: Write (Events/Clearing) - can read for read-modify-write
    // Port B: Read (Readout) - independent read port, 1-cycle latency
    // =========================================================================
    // Port A signals for write operations
    logic [CELL_ADDR_BITS-1:0] port_a_addr;
    logic [COUNTER_BITS-1:0] port_a_rdata;  // Read data from Port A
    logic [COUNTER_BITS-1:0] port_a_wdata;
    logic port_a_wen;
    
    // Port B signals for readout (read-only)
    // rd_addr is already defined above
    
    // Port A: Handle writes (clearing and events)
    // For events: Read-Modify-Write pipeline (2 cycles)
    logic event_valid_pipe;
    logic [CELL_ADDR_BITS-1:0] evt_addr_pipe;
    logic [COUNTER_BITS-1:0] evt_read_data;
    
    always_ff @(posedge clk) begin
        // Port A read (registered for read-modify-write)
        port_a_rdata <= mem[port_a_addr];
        
        // Pipeline event address and valid
        event_valid_pipe <= event_valid;
        evt_addr_pipe <= evt_addr;
        evt_read_data <= port_a_rdata;  // Capture read data for write
        
        // Port A write
        if (port_a_wen) begin
            mem[port_a_addr] <= port_a_wdata;
        end
    end
    
    // Port B: Read port for readout (independent, no conflicts)
    always_ff @(posedge clk) begin
        if (readout_busy) begin
            ram_rdata <= mem[rd_addr];  // Port B read
        end
    end
    
    // Port A address and write control
    always_comb begin
        port_a_addr = '0;
        port_a_wdata = '0;
        port_a_wen = 1'b0;
        
        if (state == S_CLEAR) begin
            // Priority: Clearing (direct write, no read needed)
            port_a_addr = clear_addr;
            port_a_wdata = '0;
            port_a_wen = 1'b1;
        end else if (event_valid_pipe) begin
            // Event Integration: Write using pipelined read data
            port_a_addr = evt_addr_pipe;
            if (evt_read_data != {COUNTER_BITS{1'b1}}) begin
                port_a_wdata = evt_read_data + 1'b1;  // Increment
            end else begin
                port_a_wdata = evt_read_data;  // Saturate
            end
            port_a_wen = 1'b1;
        end else if (event_valid) begin
            // First cycle: initiate read (address set, write disabled)
            port_a_addr = evt_addr;
            port_a_wen = 1'b0;  // Read only
        end
    end
    
    // Note on Latency:
    // `readout_valid` needs to match `ram_rdata` timing.
    // In `always_ff`, `ram_rdata` updates 1 cycle after address change.
    // `readout_busy` logic updates `rd_cell_ctr`.
    // The `ram_rdata` corresponds to `rd_addr` from PREVIOUS cycle.
    // So `readout_valid` should be delayed by 1 cycle relative to `readout_busy` start?
    // In strict pipelining:
    // Cycle 0: trigger set.
    // Cycle 1: busy=1, addr=0.
    // Cycle 2: data=mem[0] ready. valid should be 1.
    // My FSM sets `readout_valid <= 1` immediately when busy is true.
    // So on Cycle 1 (if triggered prev), valid=1. But data isn't ready.
    // I need to delay valid by 1 cycle relative to address application.
    
    logic readout_valid_d;
    always_ff @(posedge clk) begin
        readout_valid_d <= (readout_busy); // Valid if we were busy reading last cycle
    end
    assign readout_valid = readout_valid_d;

endmodule
